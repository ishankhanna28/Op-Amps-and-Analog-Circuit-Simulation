* C:\Users\Ishan's PC\Desktop\Sem 4\Lab\LIC\Differentiator\sch.sch

* Schematics Version 9.2
* Thu Mar 18 00:09:22 2021



** Analysis setup **
.tran 0ns 100
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "sch.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
