* C:\Users\Ishan's PC\Desktop\Sem 4\Schematic1.sch

* Schematics Version 9.2
* Thu Mar 11 02:28:18 2021



** Analysis setup **
.tran 0ns 5ms
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
