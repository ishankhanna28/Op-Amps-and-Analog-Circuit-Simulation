* C:\Users\Ishan's PC\Desktop\Sem 4\Lab\LIC\Integrator Practical\integratore_reale_transient.sch

* Schematics Version 9.2
* Thu Mar 18 01:14:20 2021



** Analysis setup **
.tran 0.1ms 100ms 50ms
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "integratore_reale_transient.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
